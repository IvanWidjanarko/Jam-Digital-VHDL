LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

ENTITY JAM_DIGITAL IS
	PORT
	(
		RESET				:	INOUT	STD_LOGIC	:= '0';
		CLOCK				:	IN		STD_LOGIC;
																								-- JAM = 07 (21/3)
		JAM_1				:	INOUT	STD_LOGIC_VECTOR (1 DOWNTO 0)	:=	"00";		--0
		JAM_2				:	INOUT	STD_LOGIC_VECTOR (3 DOWNTO 0)	:= "0111";	--7
																								-- MENIT = 12 roundup(23/2)
		MENIT_1			:	INOUT	STD_LOGIC_VECTOR (2 DOWNTO 0)	:= "001";	--1
		MENIT_2			:	INOUT	STD_LOGIC_VECTOR (3 DOWNTO 0) := "0010";	--2
																								-- DETIK = 36 (6*6)
		DETIK_1			:	INOUT	STD_LOGIC_VECTOR (2 DOWNTO 0)	:=	"011";	--3
		DETIK_2			:	INOUT	STD_LOGIC_VECTOR (3 DOWNTO 0)	:=	"0110";	--6
		SEVEN_JAM_1		:	OUT	STD_LOGIC_VECTOR (6 DOWNTO 0);
		SEVEN_JAM_2		:	OUT	STD_LOGIC_VECTOR (6 DOWNTO 0);
		SEVEN_MENIT_1	:	OUT 	STD_LOGIC_VECTOR (6 DOWNTO 0);
		SEVEN_MENIT_2	:	OUT	STD_LOGIC_VECTOR (6 DOWNTO 0);
		SEVEN_DETIK_1	:	OUT	STD_LOGIC_VECTOR (6 DOWNTO 0);
		SEVEN_DETIK_2	:	OUT 	STD_LOGIC_VECTOR (6 DOWNTO 0)
	);
END JAM_DIGITAL;

ARCHITECTURE DIGITAL_CLOCK OF JAM_DIGITAL IS
BEGIN

	WAKTU : PROCESS (RESET,CLOCK,JAM_1,JAM_2,MENIT_1,MENIT_2,DETIK_1,DETIK_2)
	BEGIN
		IF (RESET = '1') THEN
			JAM_1		<=	"00";
			JAM_2		<=	"0000";
			MENIT_1	<=	"000";
			MENIT_2	<=	"0000";
			DETIK_1	<=	"000";
			DETIK_2	<=	"0000";
			RESET		<=	'0';

		ELSIF(RISING_EDGE(CLOCK))THEN
			DETIK_2	<=	DETIK_2 + 1;
		END IF;

		
		IF (DETIK_2 = "1010") THEN
			DETIK_2	<=	"0000";
			DETIK_1	<=	DETIK_1 + 1;	
		ELSIF (MENIT_2 = "1010") THEN
			MENIT_2	<=	"0000";
			MENIT_1	<=	MENIT_1 + 1;
		ELSIF (JAM_2 = "1010") THEN
			JAM_2		<= "0000";
			JAM_1		<=	JAM_1 + 1;
		END IF;
		
		
		IF (DETIK_1 = "110") THEN
			DETIK_1	<=	"000";
			MENIT_2	<=	MENIT_2 + 1;
		ELSIF (MENIT_1 = "110") THEN
			MENIT_1	<= "000";
			JAM_2		<=	JAM_2  + 1;
		ELSIF (JAM_1 = "10") THEN
			IF (JAM_2 = "0100") THEN
				RESET	<=	'1';
			END IF;
		END IF;
	
	END PROCESS WAKTU;

	SEVEN_HOUR_1 : PROCESS (JAM_1) IS
	BEGIN
		CASE JAM_1 IS
			WHEN "00"	=> SEVEN_JAM_1 <= "1111110"; --0
			WHEN "01"	=> SEVEN_JAM_1 <= "0110000"; --1
			WHEN "10"	=> SEVEN_JAM_1 <= "1101101"; --2
			WHEN OTHERS	=> SEVEN_JAM_1 <= "0000000"; --TIDAK ADA
		END CASE;
	END PROCESS SEVEN_HOUR_1;
	
	SEVEN_HOUR_2 : PROCESS (JAM_2) IS
	BEGIN
		CASE JAM_2 IS
			WHEN "0000" => SEVEN_JAM_2 <= "1111110"; --0
			WHEN "0001" => SEVEN_JAM_2 <= "0110000"; --1
			WHEN "0010" => SEVEN_JAM_2 <= "1101101"; --2
			WHEN "0011" => SEVEN_JAM_2 <= "1111001"; --3
			WHEN "0100" => SEVEN_JAM_2 <= "0110011"; --4
			WHEN "0101" => SEVEN_JAM_2 <= "1011011"; --5
			WHEN "0110" => SEVEN_JAM_2 <= "1011111"; --6
			WHEN "0111" => SEVEN_JAM_2 <= "1110000"; --7
			WHEN "1000" => SEVEN_JAM_2 <= "1111111"; --8
			WHEN "1001" => SEVEN_JAM_2 <= "1110011"; --9
			WHEN OTHERS => SEVEN_JAM_2 <= "0000000"; --TIDAK ADA
		END CASE;
	END PROCESS SEVEN_HOUR_2;
	
	SEVEN_MINUTE_1 : PROCESS (MENIT_1) IS
	BEGIN
		CASE MENIT_1 IS
			WHEN "000"	=> SEVEN_MENIT_1 <= "1111110"; --0
			WHEN "001"	=> SEVEN_MENIT_1 <= "0110000"; --1
			WHEN "010"	=> SEVEN_MENIT_1 <= "1101101"; --2
			WHEN "011"	=> SEVEN_MENIT_1 <= "1111001"; --3
			WHEN "100"	=> SEVEN_MENIT_1 <= "0110011"; --4
			WHEN "101"	=> SEVEN_MENIT_1 <= "1011011"; --5
			WHEN OTHERS	=> SEVEN_MENIT_1 <= "0000000"; --TIDAK ADA
		END CASE;
	END PROCESS SEVEN_MINUTE_1;

	SEVEN_MINUTE_2 : PROCESS (MENIT_2) IS
	BEGIN
		CASE MENIT_2 IS
			WHEN "0000" => SEVEN_MENIT_2 <= "1111110"; --0
			WHEN "0001" => SEVEN_MENIT_2 <= "0110000"; --1
			WHEN "0010" => SEVEN_MENIT_2 <= "1101101"; --2
			WHEN "0011" => SEVEN_MENIT_2 <= "1111001"; --3
			WHEN "0100" => SEVEN_MENIT_2 <= "0110011"; --4
			WHEN "0101" => SEVEN_MENIT_2 <= "1011011"; --5
			WHEN "0110" => SEVEN_MENIT_2 <= "1011111"; --6
			WHEN "0111" => SEVEN_MENIT_2 <= "1110000"; --7
			WHEN "1000" => SEVEN_MENIT_2 <= "1111111"; --8
			WHEN "1001" => SEVEN_MENIT_2 <= "1110011"; --9
			WHEN OTHERS => SEVEN_MENIT_2 <= "0000000"; --TIDAK ADA
		END CASE;
	END PROCESS SEVEN_MINUTE_2;

	SEVEN_SECOND_1 : PROCESS (DETIK_1) IS
	BEGIN
		CASE DETIK_1 IS
			WHEN "000"	=> SEVEN_DETIK_1 <= "1111110"; --0
			WHEN "001"	=> SEVEN_DETIK_1 <= "0110000"; --1
			WHEN "010"	=> SEVEN_DETIK_1 <= "1101101"; --2
			WHEN "011"	=> SEVEN_DETIK_1 <= "1111001"; --3
			WHEN "100"	=> SEVEN_DETIK_1 <= "0110011"; --4
			WHEN "101"	=> SEVEN_DETIK_1 <= "1011011"; --5
			WHEN OTHERS	=> SEVEN_DETIK_1 <= "0000000"; --TIDAK ADA
		END CASE;
	END PROCESS SEVEN_SECOND_1;

	SEVEN_SECOND_2 : PROCESS (DETIK_2) IS
	BEGIN
		CASE DETIK_2 IS
			WHEN "0000" => SEVEN_DETIK_2 <= "1111110"; --0
			WHEN "0001" => SEVEN_DETIK_2 <= "0110000"; --1
			WHEN "0010" => SEVEN_DETIK_2 <= "1101101"; --2
			WHEN "0011" => SEVEN_DETIK_2 <= "1111001"; --3
			WHEN "0100" => SEVEN_DETIK_2 <= "0110011"; --4
			WHEN "0101" => SEVEN_DETIK_2 <= "1011011"; --5
			WHEN "0110" => SEVEN_DETIK_2 <= "1011111"; --6
			WHEN "0111" => SEVEN_DETIK_2 <= "1110000"; --7
			WHEN "1000" => SEVEN_DETIK_2 <= "1111111"; --8
			WHEN "1001" => SEVEN_DETIK_2 <= "1110011"; --9
			WHEN OTHERS => SEVEN_DETIK_2 <= "0000000"; --TIDAK ADA
		END CASE;
	END PROCESS SEVEN_SECOND_2;
	
END DIGITAL_CLOCK;